module qc_top(
    input  logic clk,
    input  logic start,
    output logic done
);
    scheduler sched(.clk(clk), .start(start), .done(done));
endmodule
